module contract

pub enum TypeGenerate {
	v
	csharp
}
