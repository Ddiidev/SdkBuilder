module main

import builder_sdk

fn main() {
	builder_sdk.construct(r'C:\Users\AndreLuiz\Documents\SourceApps\Vlang\SdkTest\sdkbuilder.json')!
}
